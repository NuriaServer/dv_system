`include "base_test.sv"

`include "seq_i2c.sv"

`include "test_dummy.sv"

`include "test_i2c_read.sv"