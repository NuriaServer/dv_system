`include "base_test.sv"

`include "seq_i2c.sv"

`include "test_dummy.sv"